// this is the equivalent to bigman from lab10
module isqrt (
    input [7:0] a,
    input [3:0] sqrt
);
    
endmodule