module bin2bcd (
    input [7:0] bin,
    output reg [11:0] bcd
);

//TODO: Do the thing
endmodule
