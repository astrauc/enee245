module isqrt (
    input [11:0] a,
    input clk, 
    input clr, 
    input en_a,
    input en_del,
    input en_sqrt,
    input en_out, 
    input ld_add,
    output reg [3:0] sqrt.
    output reg greater
);

    
    
endmodule