module controller (
    input greater,
    input start, 
    input clk,
    input clr, 
    output en_a,
    output en_del,
    output en_sqrt,
    output en_out, 
    output ld_add,
);


    
endmodule