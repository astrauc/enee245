module vendingMachine (

);

// Next state logic block
// This computes:
// What state do we need to go to given the current state and the inputs

// State memory block
// This computes: 
// 

// Output state logic block

endmodule